module tb;
  initial begin
    $display("Hi");
  end
endmodule
