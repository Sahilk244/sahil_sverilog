module tb;
  initial begin
    $display("I am sahil brother");
  end
endmodule
